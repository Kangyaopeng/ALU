../uvc/op_s_agent/op_s_if.sv