/***********************************************
#
#      Filename:    inst.v
#
#        Author:  Kang Yaopeng   -- 78490223@qq.com
#   Description:  ---
#        Create:  2019-03-12 15:08:20
# Last Modified:  2019-03-12 15:08:20
***********************************************/
`timescale 1ns/1ps
module inst(output out1, output out2);
  assign out1 = 1'b1;
  assign out2 = 1'b1;
endmodule
