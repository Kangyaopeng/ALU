../uvc/apb_agent/apb_if.sv