../uvc/op_m_agent/op_m_if.sv